module coffee_brewer (
    input 
);
    
endmodule