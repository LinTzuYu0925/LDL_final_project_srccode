module state_FSM (
    input clk,
    input rst
);
    
endmodule

module mode_FSM (
    input clk,
    input rst
);
    
endmodule

module water_FSM (
    input clk,
    input rst
);
    
endmodule